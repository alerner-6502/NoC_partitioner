module noc_0 (
	input  i_rst,
	input  i_clk,
	
	//connections to SUBNOC #1
	input  [7:0] i_valids_1,
	input  [7:0] i_credits_1,
	input  [7:0] i_flits_1 [7:0],
	output [7:0] o_valids_1,
	output [7:0] o_credits_1,
	output [7:0] o_flits_1 [7:0]
);

	//USER CODE FOR SUBNOC #0

endmodule

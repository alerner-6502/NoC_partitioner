module noc_1 (
	input  i_rst,
	input  i_clk,
	
	//connections to SUBNOC #0
	input  [7:0] i_valids_0,
	input  [7:0] i_credits_0,
	input  [7:0] i_flits_0 [7:0],
	output [7:0] o_valids_0,
	output [7:0] o_credits_0,
	output [7:0] o_flits_0 [7:0]
);

	//USER CODE FOR SUBNOC #1

endmodule
